-- NUT0..2.ROM

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM41C is
   port(
      OutClock      : in std_logic;
      OutClockEn    : in std_logic;
      Reset         : in std_logic;
      Address       : in std_logic_vector(13 downto 0);
      Q             : out std_logic_vector(9 downto 0)
   );
end ROM41C;

architecture logic of ROM41C is
    type mem_t is array(0 to 16383) of integer range 0 to 1023;
    constant rom : mem_t := (
      
         513,    6,  693,    6,   78,  624,  248,  344,  920,   86,  644,  984,  332,   91,  140,   75, 
          76,   59,  796,   66,  624,  112,   56,   75,  174,  888,   60,  518,  112,  441,   88,  206, 
         652,  928,  909,    8,  644,  923,  630,  630,  537,    8,  174,  856,  764,   88,  243,  409, 
         158,  665,   10,  693,  150,  269,  158,   21,  150,  189,  150,  610,  610,  966,  970,  592, 
          28,   35,  537,    8,  174,  856,  764,   88,  482,   27,  482,  311,   17,    0,  238,  860, 
         152,   28,  581,    2,  652,  928,  644,   17,    0,  909,    8,  856,  268,  928,  181,  162, 
         635,  155,  715,  707,  275,  227,  219,  331,  323,  715,  571,  579,  587,  595,  603,  701, 
         178,  337,    0,  739,  270,  540,  848,  790,  693,   35,   17,   12,  174,  270,  147,  964, 
         131,  112,  506,  368,  672,   51,  240,  184,  270,  865,   80,  248,  869,   80,  964,  240, 
         124,  304,   20,  636,  816,   80,  444,  480,  968,  972, 1015,  304,    8,  968,  972,  614, 
        1003,  992,  981,  136,   79,  165,   80,  240,  212,   79,  165,   80,  212,   63,  168,  240, 
         238,  459,  165,   80,  174,  952,  380,  856,  174,  652,  935,  332,  819,  324,  920,  316, 
         936,  387,  949,  444,  388,  355,  588,  609,    0,  323,   19,    0,  165,   80,  238,  212, 
         211,  952,  380,  856,  652,  819,  163,  432,  368,  992,  165,   80,  238,  212,   51,  952, 
         380,  856,  652,  707,  120,  168,   78,  624,   56,  104,  248,  296,  238,  232,  949,  444, 
         392,  608,  160,   78,  624,  952,  856,  352,   67,  332,   55,  328,  237,    4,  369,   28, 
         748,   31,  524,   27,  913,  156,  716,  411,  972,  163,  544,   60,   86,  262,  304,   24, 
         870,  801,   70,  304,  135,  870,   47,  529,   12,  797,    2,  968,  972,   92,   90,  976, 
         368,  824,  204,  151,  260,  610,   71,  808,  624,  124,  304,   20,  252,  480,  400,  614, 
         808,   28,  624,   56,  283,  558,  808,  444,  816,  235,  307,  952,  920,  936,  992,    0, 
         163,  131,   99,   67,   35,   56,  892,  131,   56,  252,  107,   56,  316,   83,   56,  380, 
          59,   56,  124,   35,   56,  264,  572,  908,   27,  941,  444,  304,    6,  624,  252,  480, 
         584,  369,   28,  140,  127,   12,   35,  393,   20,   83,  652,   43,  260,   65,  176,   35, 
         248,  153,   44,  588,   63,  304,   81,  614, 1019,  609,    0,   68,  237,    4,  780,  199, 
           1,  256,  981,   12,  972,  271,  304,    8,  921,  156,  524,  975,  952,  572,  856,   12, 
         985,   28,   96,    0,  369,   28,  747,  345,   36,  304,   92,  262,  972,   79,  304,   12, 
         945,  156,  422,  971,  777,   30,  544,   28,  482,   21,   50,  801,   70,    1,  256,  736, 
         981,   12,  972,   63,  304,   10,  921,  156,  524,  699,  952, 1009,   12,  380,  984,  772, 
         136,  324,  644,  984,  572,   70,  380,  936,  708,  888,  238,  304,  191,  270,  358,  806, 
         123,  166,  262,  624,   56,  750,   75,  574,  951,   94,  752,  252,   86,  326,  907,  304, 
           7,  624,  921,  156,   81,  132,   78,  624,  609,    0,  972,   75,  304,  195,  262,  544, 
          60,  796,  874,  507,  800,  952,  444,  856,  908,  965,    2,  900,  920,   60,  936,  736, 
         877,   88,  800,  777,   30,  968,  972,  608,   70, 1008,  624,  304,  361,  262,  888,  380, 
         870,  271,  444,  614,  624,   56,  270,  698,  752,   56,  698,  878,  183,  752,   70,  624, 
         952,  856,  204,  928,  824,   70,  444,  816,  742,  864,  196,  888,   60,   28,   66,  266, 
         189,  142,  608,  416,  344,  112,   88,  856,  600,  368,  368,  368,  368,  224,  732,  160, 
         708,  836,  388,  196,  580,  260,  433,  112,   45,  985,   28,  609,    0,  304, 1023,  270, 
          78,  752,  736,  800, 1008,  174,  624,  174,  752,  422,  987,  304,  239,  316,  304,  250, 
          60,  304,  238,  872,   90,  558,  808,  624,   78,  156,  784,  304,   32,  936,   78,  624, 
         668,  144,  784,   92,  272,  528,  936,  136,  304,    6,  921,  156,  304,  361,  262,  888, 
         380,  166,  316,  872,  981,    6,  270,  716,   31,   76,  928,  824,  204,   67,  558,  808, 
         444,  816,  182,  262,  992,  268,  107,  400,  614,  808,  624,   56,  892,  796,  266,   28, 
          78,  624,  992,  610,  808,  992,  537,    8,  174,  856,  540,   88,  502,  701,  190,  580, 
         502,   67,  584,  502,   43,  502,  864,  317,    2,   86,  652,   51,  644,   17,    0,  945, 
          14,  174,  142,  304,   30,  454,   63,  588,  195,  304,   26,  454,  163,  110,  304,    8, 
         238,   78,  624,  558,  572,  390, 1011,   19,  494,  358, 1011,  238,  952,  174,  317,    2, 
         981,  136,   56,  638,  638,  905,   83,  262,   94,  260,   70,  624,  854,  864,  892,  422, 
          71,  264,  764,  422,   39,  764,  422,  843,  572, 1005,    8,  486,  262,  486,  486,  326, 
          70,  764,  518,  992,   28,  142,  206,  716,   71,   76,   55,  632,  588,   23,  344,  992, 
         204,  387,  824,  444,  570,  238,  482,  223,  206,  816,  142,  282,  828,  638,  286,   78, 
         796,  174,  570,  816,  174,  170,  572,  446,  971,   19,  572,  746, 1011,  344,  174,  110, 
          28,   83,  206,  570,  816,  828,   70,  252,  110,  538,  570,   60,  234,  824,  202,  808, 
         992,  580,  482,   51,  329,  164,  857,  164,   27,  329,  164,  741,  164,  828,  286,   78, 
         446,   79,  344,  741,  164,  984,  408,  984,  572,  955,  805,   80,  344,   28,  221,  140, 
         110,  952,  856,  992,  869,  444,  652,   27,  716,  928,  260,  584,   65,  176,   51,  877, 
         444,  206,  153,   44,  505,   12,  908,   47,  316,  856,  524,  359,  613,   32,   70,  624, 
         952,  856,  136,  211,  708,  952,  572,  856,  772,  920,  892,  856,  772,   43,  329,   36, 
         952,  856,  380,  984,  772,  984,  252,  984,  900,  516,  984,  892,  132,  920,  936,  992, 
         901,  444,  569,   12,  260,  652,  443,  952,  856,  772,  237,    4,  708,  992,  432,  538, 
         816,  742,  283,   28,   80,  444,  174,  961,  176,  174,  845,   20,  989,  172,  329,   36, 
         613,   32,  861,  444,  357,   28,   76,  629,   46,  952,  856,  136,  920,  380,  856,  776, 
         920,  316,  936,  797,    2,  952,  856,  132,  920,  380,  856,  772,  931,   65,  176,  505, 
          12,  563,  304,  167,  968,  972,  761,   30,  614,  987,  557,  170,  909,    8,  758,  897, 
          11,  540,  152,  689,   10,  304,  765,  624, 1008,  184,   21,   10,   70,  936,  777,  186, 
         139,  163,  171,  219,  179,  171,  163,  155,  147,  251,  419,  243,  259,  299,  291,  969, 
          18,  304,  207,  422,   99,  693,   18,  304,  144,   59,  797,   20,  521,   18,  304,  145, 
           2,  134,  262,  797,   20,  102,  900,  483,  371,  304,  208,  835,  304,  206,  774,  355, 
         101,   22,  924,    2,  797,   20,   17,  180,   29,  180,  984,  644,  984,  283,  304,  168, 
         774,  297,  191,  304,  174,  774,  175,   25,  180,  984,  985,   28,  652,   35,  304,  224, 
          27,  304,  208,  813,   20,  147,  904,  304,  156,  774,   19,  900,  797,   20,   17,  180, 
         262,  985,   28,  166,  984,  652,  115,  644,  984,  900,  230,  957,   28,    9,   14,  516, 
         733,   20,  102,   27,  984,  262,   22,  304,  102,  774,  107,   30,  382,  908,   23,  382, 
         929,   20,  780,  989,  172,  605,   30,  304,  112,  774,  199,  870,  139,  304,  116,  870, 
         211,  774,  155,  304,  113,  582,  828,  304,   26,  638,   55,  614, 1003,  304,   92,  582, 
        1000,  779,  304,  101,  987,  304,  122,  582,  566,  955,  304,  104,  923,  304,   29,  774, 
         459,  315,  304,   26,  774,  207,  870,  103,  952,  984,  328,  348,  162,  482,   23,  648, 
         984, 1000,  139,  550,  870,   55,  733,   20,  304,    5,   59,  304,   45,   35,  166,  796, 
         208,  741,   20,   17,  180,  110,   86,  262,  985,   28,  304,   29,  796,  866,   31,  774, 
         663,  268,   43,  304,   31,  741,   20,  521,   18,  998,   22,  797,   20,   17,  180,  110, 
         262,  260,  516,  204,   19,  520,  796,    2,  166,   90,   86,  444,  282,  985,   28,  952, 
         304,  263, 1000,  442,  751,  110,  329,   36,   28,  524,   45,  181,  524,  741,  164,  110, 
         262,  985,   28,  166,  373,  176,  745,   20,  859,  110,  829,  164,   29,  180,  142,  262, 
         985,   28,  796,  354,  115,  304,  207,  813,   20,  329,   36,  110,  829,  164,  110,  430, 
         965,   18,  170,  610,  856,  304,  192,  813,   20,  204,  239,  140,  219,  736,  952,  952, 
         304,   68, 1000,  617,   20,  262,   30,  985,   28,  929,   20,  304,   32, 1000, 1016,  924, 
         738,   19,  936,  304,   96,  936,  800,  772,  339,  304,  200,  584,  968,  972,  928,  614, 
         995,  580,  260,  772,  900,  329,   36,  557,  168,  262,  134,  844,   43,  429,  112,   67, 
         147,  961,  176,   30,  929,   20,  710,  111,  204,   79,  617,   20,  262,   30,  985,   28, 
         929,   20,  521,   18,  304,   32, 1000,  329,   36,  952,  270,  321,  164,   29,  180,  796, 
         746,  995,  142,   86,  262,  572,  304,   64,  252,  480,  957,   28,   32,   18,    5,    7, 
         544,  329,   36,  888,   90,  270,   67,  614,  270,  624,   56,  750,   71,  378,  304,  192, 
         870,   27,  174,  931,  174,   60,  992,  304,   32, 1000,  780,   87,  304,   32,  262, 1016, 
         936,   86,  870,  928,  776,  889,  178,  985,   28,  166,  262,  572,  304,   20,  636,  816, 
          28,   80,  444,  264,  634,  816,   86,  984,  332,   27,  566,  324,  652,   27,  260,  644, 
         984, 1000,  268,  911,  304,   32, 1000,  992,  158,   78,  672,  166,  270,  572,  550,  614, 
         494,  494,  494,  494,  998,  166,  572,  550,  614,  518,  190,  494,  494,  494,  494,    6, 
         174,  764,  558,  622,  526,  608,  734,  119,  732,  272,  286,  124,  766,  127,  764,  446, 
         766,   95,  764,  446,   67,  126,  158,  446,   31,  828, 1003,  126,  828,  282,  158,  764, 
         924,  446,  864,  304,    3,  764, 1000,  979,   70,  624,  206,  493,   40,  260,   20,   19, 
         264,  174,  344,  766,  973,  125,  224,  860,  224,  724,  864,  208,  988,   98,  770,  215, 
         866,  147,   98, 1001,  124,  224,  194,  482,   35,  304,   44,   27,  304,   46,  980,  160, 
         981,  124,  819, 1001,  124,  224,  980,  532,  771,  268,  928,  796,  408,  738,   23,  980, 
         160,  304,   69,  981,  124,  408,  758,  973,  125,  635,   28,  824,  444,  836,   19,  634, 
         816,  630, 1007,  630,  991,  630,   23,  840,   60,  266,  992,  204,   27,  170,  883,  313, 
         136,  742,  777,   82,  213,  136,  574,  983,  845,  166,  293,   28,  985,   28,  304,   32, 
        1000,  277,   56,    0,  332,  115,  176,  482,   47,  304,   45, 1000,   19,  952,  917,  124, 
         985,   28,  891,  304,  195,  270,  544,   60,  778,   35,  613,   32,  811,   78,  544,   60, 
         208,  550, 1000,  262,  304,   52,  260,  870,   23,  264,  176,  966,  262,  966,  796,  208, 
         268,   27,  738,   23,  546, 1000,  358,  497,   58,  270,  304,   65,  774,  864,  304,   75, 
         774,  243,  304,   37,  518,  764,  230,  796,  266,  304,   30,  874,   35,  614,  874,   55, 
         252,  270,  102,  641,   58,  304,  205,  874,   47,  828,  574,  574,  931,  102,  992,  304, 
          97,  774,  864,  304,  102,  774,  928,  304,   26,  731,  176,  828,  270,  358,  772,  513, 
         172,   12,  271,   28,  738,   47,  270,   22,  657,   62,  112,    1,   32,   83,  174,  472, 
          12,   39,  176,  689,   62,  520,  395,  961,  176,  433,  188,  329,   36,  580,  176,  929, 
          28,  505,   62,  344,  925,  444,  408,   28,  285,  136,  764,  286,  446,  446,  733,  164, 
          78,  112,  741,  164,  984,  176,  984,  572,  446,  963,  805,   80,  112,   70,  624,  176, 
         616,  304,   30,  892,  929,   28,  516,  501,   62,  952,  828,  984,   68,  984,  764,  936, 
         985,   28,  376,  984,  644,  984,  752,  329,   38,  577,   12,  936,  304,  128,  166,  998, 
          78, 1008,  624,  952,  856,  716,   31,   12,   27,  358,  358,  332,   23,   22,  652,   19, 
         366,  572,  856,  908,   35,  304,  128,  326,   76,   47,  140,   35,  374,  374,  374,  188, 
         856,  908,   43,  374,  374,  374,  374,  188,   86,  494,  828,   86,  494,  494,  334,  304, 
          16,  624,  304,  253, 1008,  174,  752,   70, 1008,  624,  952,  856,  992,  380,  984,  780, 
         733,   47,  856,   12,   43,  304,  132,  589,   50,  780,  991,  905,   12,  844,   51,  260, 
         433,  112,   67,   75, 1016,  742,   31,  550, 1000,  357,   20,  588,  793,   56,  893,  444, 
         357,   28,  712, 1016,   70,  614, 1000,  952,  856,  502,  502,   43,  925,  444,  577,   12, 
         772,  952,  920,  936,  345,   36,  140,   71,  961,  176,  304,   46,  936,  329,   36,  961, 
           2,   78,  552,  488,  424,  152,  360,  992,  764,   92,  266,  696,  170,  680,  992,  432, 
         816, 1000,  570,  758,  995,  480,  304,   16,  624,  304,  253, 1008,  992,    0,    0,    0, 
          90,  494,  494,  764,  966,  486,  486,  966,   60,  262,  444,  348,  234,   90,  336,  348, 
         816,  870,   35,  546,  995,  992,  570,  198,  270,  816,  550,  774,  195,  166,  486,  378, 
          90,  444,  538,  816,  502,  502,  572,  856,  252,  270,  572,  570,  816,  796,  266,   60, 
         346,  432,  570,  480,  634,  755,  260,  568,  444,  856,  860,  152,  766,  661,   38,  764, 
         784,  720,  656,  270, 1006,  894,  403, 1006,  780,  561,   35,  894,  219, 1006,  894,  163, 
         766,   19,    8,   28,  632,  546,   27,  988, 1003,   20,  613,   35,  908,   39,  632,  638, 
         616,  641,   34,  908,  431,  904,  219,  632,  270,  732,  144,  798,  367,  776,   12,  455, 
          78,  622,   86,  732,  592,   80,    8,  379,  780,   95,  268,   31,   12,  227,  524,   31, 
         520,  307,  516,  291,  632,  270,   86,  540,  854,   23,  848,  219,  894,   99, 1006,  894, 
          75,  924,  632,  546,   27,  988, 1003,  916,   67,  736,  304,  208,  614, 1019,  800,  992, 
         980,    0,  152,  258,  632,  162,  616,  568,  444,  920,   60,  552,  992,  540,  174,   88, 
         264,   19,  260,   78,  622,   86,  732,  656,  616,  653,  184,  952,  856,   12,   43,  713, 
         140,  649,  182,  396,  949,   81,  392,   78,  232,  268,  477,  182,  321,  164,  138,  329, 
          36,  221,   32,  377,   36,   25,  180,  106,  796,  266,  304,   29,  866,   63,  778,   43, 
         174,  924,   88,  867,  110,  797,  164,  221,  140,  961,    2,  110,  608,   28,  971,  568, 
         444,  856,  632,  270,  985,   28, 1001,   80,   28,  354,   43,  610,  446,  988,  987,  418, 
         780,   71,   20,   55,  980,  418,   80,  988,  988,  908,   91,  446,   31,  988, 1003,  140, 
          27,  464,   19,  976,  988,   76,  155,  724,  127,  286,  446,   47,  852,  103,  988,  987, 
         140,   27,  976,   19,  464,  988,  923,  190,   19,  286,  446,   94,  732,  524,   19,  848, 
         190,  224,  732,  160,  630,  780,  131,  796,  354,   71,  418,  924,  354,   47,  418,  546, 
          35,   10,  418,   80,   28,  992,   22,  924,  992,  978,  978,  104,  174,  978,  978,   40, 
          78,  168,   70, 1008,  624,  992,  985,   28,  376,  984,  776,  984,  752,  939,  632,   28, 
         546,   27,  988, 1003,  610,  262,   86,  924,  354,   43,  966,  988,  532,  987,  672,  854, 
          19,  646,  270,  732,  592,  190,  478,  119,  834,  119, 1018,  446,  995,  422,  834,  111, 
         638,  263,  422, 1018,  979,   30,  955,  446,   39,  358, 1003,  995,   30,  524,   19,  446, 
         174,  780,  131,  165,   80,  232,  852,  103,  268,  941,   35,  853,  444,  577,   12,  797, 
           2,   78,  232,  608,  992,  632,  224,  860,  160,  286,  780,   27,  924,   19,   28,  546, 
          43,  610,  446,  988,  987,  780,  131,  532,   71,   66,  754,   31,  516,    4,  976,  267, 
         630,  630,   19,  772,   86,  219,  724,   95,  908,   47,  852,   63,  574,  867,  446,  851, 
         900,  131,  952,  856,   12,   43,  577,   12, 1021,  138,   78,  232,   32,  304,  119,  992, 
         616,  669,   34,  580,  376,  796,  746,  305,  182,  270,  440,  170,  174,  572,  360,  504, 
         170,  174,  572,  424,  568,  170,  174,  572,  488,  568,  380,   74,  252,  552,  632,  766, 
         315,  265,  184,  952,  984,  332,   87,  652,   71,  984,  222,  574,  254,  305,  184,  243, 
         324,  644,  984,  262,  304,   32,  870,   87,   70, 1008,  624,  568,   86,  870,   55,  985, 
          28,  166, 1000,  851,  985,   28,  803,  264,   65,  176,  206,  365,  184,  793,    2,  952, 
         572,  856,  262,  248,  260,  672,  150,  860,  532,  295,  980,  438,  995,  270,  758,  299, 
         652,   99,  988,  852,  287,  358,  995,   51,  980,  532,  335,  422,  995,   46,  138,  314, 
          91,  270,   10,  262,  796,  554,   79,   14,  382,  910,  412,   10,  186,  608,  992,  174, 
         854,  995,   70,  931,  652,  835,  795,  358,   35,  154,  314,  823,  268,   31,   78,  883, 
         644,  118,  555,  268,  843,    6,  924,  418,  774,  959,  795,  238,  608,  653,  184,  206, 
         264,  213,   40,  238, 1001,   80,  558,  270,  672,  952,  188,  238,  126,  230,  198,  766, 
          27,  732,  848,  652,  885,   42,  860,  758,   91,  117,   44,   85,   44,  980,  986,  446, 
         550,  995,  123,  614,   31,  980, 1003,   70,  446,  319,  117,   44,   85,   44,  980,  532, 
          71,  446,  995,  980,  532,   31,  418,  995,  924,  224,   76,   67,  126,  158,  446,   71, 
         988,  724,  995,  732,  160,  126,  131,  162,  140,   27,  976,   19,  464,  988,  162,  875, 
          85,   44,   76,  117,   45,  755,  446,  438,  174,  608,  238,  605,   30,  860,  332,  403, 
         262,  304,    3,  854,   47,  454, 1019,  326,  295,  326, 1019,  198,  646,  518,  422,   55, 
         980,  446,  995,   30,  979,  117,   44,  980,  532,   63,  446,  995,  418,  980,  532, 1003, 
         726,   27,  540,  848,   28,  166,  304,  819,  166,  224,  781,   42,  198,  166,  454,  166, 
         755,    6,  758,  711,  779,  224,  732,  288,   31,  980, 1003,  160,  992,  162,  140,   27, 
         464,   19,  976,  988,  162,  992,  160,   30,  382,  894,   67,  493,   40,  985,   28,  238, 
         293,   38,  732,  784,  254,  736,  732,  976,  976,  892,  112,  985,   28,  176,  892,  112, 
         262,  796,  842,  979,  362,   39,  373,  176,  939,  304,   32,  222,  638,   35,  800,  329, 
          38, 1000,  979,   78,  102,  422,  570,  348,  272,  348,  546,  853,   15,  816,  454,  987, 
         326,   26,  174,  444,  506,  538,  570,  816,  230,  570,  816,  572,  198,  796,   60,  162, 
         444,  514,  502,  502,  502,   39,  636,  729,   14,  892,  174,  520,  793,  188,  761,   14, 
         174,  856,  337,    0,   14,  568,  156,  266,  920,  828,  190,  174,  552,  568,  252,  550, 
         900,  230,  198,  124,  552,  638,  638,  359,  638,  333,   47,  525,   78,  304,  256,  238, 
         972,  123,  544,   60,   86,  262,  924,  482,  801,   71,  304,  135,  870,  805,   14,  968, 
         238,  614,  875,  723,  997,   92,  699,  609,    0,  675,  997,   92,  904,  568,  252,  614, 
         742,  647,  619,   28,  196,  230,  614,  614,   75,  777,   80,  272,  900,   28,  238,    1, 
          48,  321,  164,  888,  400,   28,  908,   71,  874,  853,   14,  845,  164,  829,  164,  157, 
         164,  908,   31,  124,  170,  177,  140,  961,  176,  772,  541,   20,  761,   14,  165,   80, 
         238,  212,   75,   70,  624,  952,  380,  856,  652,  749,    2,  176,  624,  238,  752,  992, 
          78,  744,  808,  106,  179,  952,  828,  856,  416,  544,  188,  304,  193,  252,   28,  480, 
           0,   16,   91,   80,   75,  144,   59, 1011,  208,   35,  189,  142,  272,  828,  262,   76, 
          35,  304,  128,  518,  112,  140,  387,  174,  796,  482,  494,  494,  494,  764,  348,   80, 
         816,  828,  486,  486,  270,  924, 1016,   60,   88,  322,  166,  856,  580,  985,   28,  304, 
          32,  262,  134,  796,  952,  874, 1011,  426,  874,   55,  198, 1000,  936,  952,  979, 1016, 
         382,  864,  446,  432,  570,  480,  262,  952,  856,  652,   35,  304,  341,  371,  380,  856, 
          76,  307,  517,  188,  750, 1001,   27,  952,  856,   12,  223,  176,   90,  572,  262,  304, 
         102,  638,  103,  924,  720,  766,   67,  796,  464,  574,  510,   83,  766,   71,  518,  344, 
         270,  205,  144,  750,  391,  176,  270,  952,  856,  304,  336,   94,  892,  518,  892,  816, 
         630,  177,  181,  444,  238,  696,   92,  202,   70,  680,   12,   43,  738,   27,  796,  546, 
         924,   88,  856,  206,  188,  304,   20,  636,  816,   28,   80,  444,  344,  368,  816,  742, 
         231,  952,  856,  992,  472,  166,  134,  293,   28,  961,  176,  304,  224,  813,   20,  772, 
         541,   16,  304,  224,  924,   88,  444,  270,  102,  584,  573,   58,  580,  293,   28,  797, 
          60,  408,  845,   20,  408,  634,  816,  758,  581,   58,  502,  502,  278,  634,  816,  534, 
         572,  856,    4,  984,  924,  162,  152,  162,   88,   12,  403,  289,   56,  299,   76,  849, 
          55,   12,   51,  189,   56,  613,   32,  931,  524,  437,   55,  332,  713,   55,  780,  951, 
         652,  973,   55,  908,  911,  862,  891,  304,  145,  174,  764,  924,  322,  605,   28,  174, 
         589,   50,  961,  176,  369,   28,  925,  444,  529,   12,  797,    2,  908,   27,  780,  179, 
         277,   56,  899,  908,  107,   76,  245,   59,   12,  245,   59,  332,  713,   55,  613,   32, 
         899,  140,  869,   59,  979,  301,   56,  731,   76,  833,   55,   12,   51,  897,   52,  613, 
          32,  931,  544,   60,  266,  304,  131,  874,  127,  304,   49, 1000,  301,   56,   59,   12, 
         897,   53,  613,   32,  963,  952,  763,  780,  827,  652,  103,  140,  795,  329,   36,    6, 
         422,  422,  696,  166,  680,  259,  952, 1016, 1000,    6,  422,  497,   59,  329,   36,  696, 
          60,  270,  908,  167,  304,  205,  140,   47,  985,   28,  981,   50,  170,  174,  444,  680, 
         152,  856,  136,  920,   88,  869,   58,  332,   83,  304,  174,  170,  174,  444,  680,  780, 
         343,  283,  304,   30,  780,  779,  614,  652,  755,  924,  152,  984,   68,  984,   88,  796, 
         304,    1,  170,  174,  444,  680,  961,  176,  304,  208,  813,   20,  936,  304,   96, 1000, 
         213,   54,  329,   36,  924,  152,  984,  328,  984,   88,  985,   28,  957,   28,    9,   14, 
           4,  544,  289,   56,  363,   76,  119,  652,  351,   12,   27,  189,   56,  613,   32,  923, 
         304,   48, 1000,   27,  304,   48,  862,   23,  558, 1000,  828,  190,  764, 1000,  405,   58, 
         190,  764,  208,   86, 1000,  289,   56,   67,   12,   27,  189,   56,  613,   32,  955,  952, 
         992,   73,   54,  957,   28,   19,   20,  544,  277,   56,  955,  304,   32,  936,  936,  936, 
         877,  124,  732,  272,  270,  304,   76,  870,  207,  545,  176,  989,  172,  329,   36,  924, 
         152,  856,  696,  540,  464,  332,   27,  540,  976,  174,  892,  162,  641,   58,  613,   32, 
         667,  304,   87,  446,  862,   43,  550,  870,  991,  771,  304,   84,  870,  739,  899,   78, 
         190,  764,  796,  208, 1000,  277,   56,   99,   12,   39,  613,   32,  971,   78,  190,  764, 
         208, 1000,  283,  952,  992,  304,   31,   67,  304,   31,   35,  304,   31, 1000, 1000, 1000, 
         989,  172,  329,   36, 1016,   28,  152, 1000,  952,  828,  856,  136,  776,  920,  764,  365, 
          28,  609,    0,  529,    6,  732,  976,  796,  270,  952,  382,  856,   76,  999,    6, 1016, 
          66,   86,  326,  446,   71,  166,  486,  262,  486,  486,  326,  931,  924,  152,  856,  332, 
          35,  304,  128,  326,  134,  989,  172,  329,   36,  696,  270,  140,  167,  102,  134,  998, 
         131,  989,  172,  329,   36,  696,  270,  304,  200,  736,  968,  972,   59,  614,  995,  800, 
         793,   56,   67,  621,    0,  961,  176,  800,  329,   36,  917,  444,  529,   12,  924,  152, 
         984,   76,   59,  844,  287,  174,  188,  977,  166,  984,   78,   92,  976,  368,  174,  188, 
         766,  365,    7,  102,  581,    2,  304,  576,  486,  968,  972,  621,    2,  614,  987,  260, 
         433,  112,   60,  304, 1000,  614, 1019,   89,   54,  329,   36,  933,  444,  952,  984,  648, 
         984,  936,   78,  616,  985,   28,  277,   56,  115,  332,  209,   62,  917,  124,  947,  605, 
          28,  644,  920,  936,   73,   54,  329,   36,  632,  750,  939,  892,   74,  616,  293,   28, 
         985,   28,  952,  795,  780,  459,  613,   32,  739,  877,  124,  262,  293,   28,  438,  955, 
         796,  304,  127,  874,  915,  304,   58,  874,  883,  304,   46,  874,  851,  304,   44,  874, 
         819,  632,  746,  799,  170,  266,  572,  616,  238,  985,   28,  545,  176,  691,    0,    0, 
           0,    0,    0,    0,  329,   36,  140,  659,  796,  632,  750,  587,  805,   80,  616,  952, 
         856,  644,  920,  365,   28,  696,   60,  262,  304,   15,  874,  553,   26,  134,  985,   28, 
         989,  172,  329,   36,  632,  224,  732,  160,  540,  754,  805,   24,  102,  304,   30,  796, 
         874,  463,  632,  344,  789,  152,  750,  143,  952,  856, 1016,   60,  924,   88,   12,  351, 
         696,  270,  917,  444,  529,   12,  897,   10,  588,  311,  344,  124,  112,  584,  132,  524, 
          43,  136,  176,  929,   28,   68,  952,  984,   12,   35,  856,   72,  920,  856,  924,   88, 
         588,   75,  797,   60,  329,   36,  408,  270,  797,  188,  696,  270,  134,  641,   58,  140, 
          83,  124,   86,  270,  952,  856,  174,  580,  589,   50,  344,  124,  929,   28,  952,  856, 
         796,  408,  444,  344,   12,   91,  816,  742,   27,  208,   59,  570,  816,  742,   23,  480, 
         144,   16,  856,  924,   88,  821,   50, 1016,  230,  961,  176,   76,  928,  102,  358,  844, 
          19,    6,   30,  929,   20,  304,   32, 1000,  992,  608,  432,  816,   51,  608,  432,  816, 
         570,  368,  494,  494,  986,  986,  986,  494,  494,  892,  480,  321,  164,  344,  845,  164, 
         749,  164,  984,  992,  860,  248,   74,  270,  446,  446,   23,   80,  817,    2,    7,  294, 
        
          65,   70,  256,    0,    2,    1,    3,    4,   66,   71,    0,    0,   39,   36,   33,   32, 
          67,   72,    0,    0,   40,   37,   34,  512,   68,   73,    0,    0,   41,   38,   35,    0, 
          69,   64,    0,   15,  128,    0,    0,  152,   30,   25,  176,   69,  108,  355,  171,   19, 
          13,    8,  176,  713,  100,  240,  184,  713,  100,  270,  176,   29,   96,  136,  713,  100, 
         203,  173,   19,   13,    8,  176,  702,  240,  851,  171,  176,   99,  132,   15,   13,  176, 
         369,  100,   59,  173,  176,  702,    0,   29,   96,  873,    2,  170,  176,  309,   96,  979, 
         165,  422,  422,  176,  309,   96,  817,    2,  178,   30,   24,  176,  270,  955,  175,  176, 
         609,   96,  827,  147,    2,    1,  176,   94,  992,  147,   15,    3,    1,  849,  132,  904, 
         776,  520,  513,  118,    0,  644,  565,  146,  140,    3,  274,  513,  601,   90,  134,    8, 
          19,    1,  289,   94,  142,    9,   19,    1,  849,  132,  819,  142,   19,  257,  425,  158, 
         143,   20,  275,  513,  369,   94,  142,    1,   20,    1,  849,  132,  683,  151,    5,    9, 
          22,    1,  401,   14,    0,  648,  643,  144,    5,    5,    2,  304,    7,  837,   90,  148, 
          19,    2,    0,  321,  138,  148,  769,  259,  513,   46,  646,  515,  309,   90,  129,   12, 
           3,   78,  360,  424,  488,  552,  992,  143,   20,  531,  408,  752,  992,  132,   12,    3, 
         577,   12,  849,   30,  144,   12,  259,  561,  138,  135,   18,   12,    3,  264,  205,   94, 
         206,   12,    3,  705,   82,  148,   19,   12,    3,   78,   40,  104,  168,   43,  152,   12, 
           3,   78,  232,  777,    2,  153,   16,   15,  259,  405,  134,  146,   45,    4,  176,  517, 
         102,  135,    5,    4,  113,   94,  132,    1,   18,    7,  153,   94,  132,    1,   18,  137, 
          94,  140,  261,  260,  673,  138,    0,    0,  701,  138,  133,  275,  516,  637,   86,  132, 
          14,    5,  135,  782,  261,  328,  769,   90,  158,   18,    5,   20,   14,    5,  949,   80, 
         184,  232,  785,    2,  152,   30,    5,  176,   41,  106,  150,    4,    1,  885,  444,  992, 
         148,    3,    1,    6,  176,  945,   98,  191,  515,  518,  174,  686,  174,  299,  177,   45, 
          24,   30,    5,   72,  176,   41,  106,  131,   63,  515,  518,  309,   88,  875,  152,  777, 
         262,  648,  769,   90,  148,   14,    9,  136,   35,  131,   18,    6,  176,  237,  102,  191, 
         531,  518,  277,   90,  131,   63,  531,  518,  309,   88,  963,    0,  357,  166,  143,  788, 
         775,  146,    8,  176,  713,  102,  147,   13,    8,  136,  971,  135,  275,  521,  900,  641, 
          86,  140,    2,  780,  142,   12,  176,  277,  110,  135,   15,   12,  136,  971,  150,    5, 
           4,   19,   65,  116,   59,  142,    1,    5,   13, 1017,  112,  661,    2,  144,   45,   18, 
         849,  132,  293,  116,  955,  134,    6,   15,  736,  304,    9,  921,  156,   21,    8,  609, 
           0,  577,    6,  152,   47,   49,  176,  557,   98,  146,   45,   16,  849,  132,  776,  520, 
         469,  120,  715,  139,    3,    1,   16,    1,  130,  136,    3,   37,  190,  702,  190,  176, 
          29,   96,  358,  358,  184,  617,   96,  817,    2,  133,   19,   16,  716,   35,  776,  237, 
           4,  689,   14,  148,   16,   13,   15,   18,   16,  641,   14,  132,   45,   18,  176,  561, 
         102,  144,   15,   20,   19,  677,   14,    0,    0,  629,   30,  152,   43,   49,   14,   12, 
         176,  461,  110,  152,   20,   19,    1,   12,  312,  238,   35,  140,  259,  530,  396,  949, 
          81,   78,  624,  238,  232,  953,    2,  147,    8,    3,  176,  762,   27,  702,  232,  947, 
         137,   16,  672,  617,  100,  494,  570,   70,  779,  190,  316,  536,  408,  752,  795,  142, 
           4,   18,  757,   82,  132,   14,   18,  189,   42,  142,   20,   18,   13,  158,  158,   18, 
         917,   82,  137,  771,  275,  769,   90,  646,  531,  297,   90,  171,   78,  545,  114,  173, 
          78,  136,  987,  135,    5,  530,  590,  357,   90,  147,   15,    3,  849,  132,  107,  142, 
           1,   20,  849,  132,   67,  142,    9,   19,  849,  132,  904,  776,  481,  122,  133,   26, 
         265,  275,  597,   94,  148,   18,   17,   19,  176,  761,   98,  148,   19,   19,    0,  385, 
         138,  142,   15,   69,   82,  170,  276,  531,  841,   80,  309,   96,   67,  171,  276,  531, 
         841,   80,   29,   96,  953,   46,  173,  276,  531,  408,  672,  702,  344,  923,  175,  276, 
         531,  841,   80,  609,   96,  891,  152,   30,   48,   49,  993,  110,  133,   14,  783,  276, 
         889,   90,  151,    5,  265,  534,  445,   14,  191,   48,   77,   24,   69,   90,  191,   25, 
          77,   24,  165,   90,  191,   48,   60,   24, 1001,   86,  191,   48,   61,   60,   24,   37, 
          90,  191,   25,   61,   60,   24,    5,   90,  153,   62,   60,   24,  248,  174,  184,  232, 
         174,  168,  953,    2,  191,   25,   60,   24,  957,   86,  191,   48,   61,   24,   25,   90, 
         191,   25,   61,   24,   81,   90,  191,   48,   62,   24,  965,   86,  191,   25,   62,   24, 
         993,   86,    0,  797,  146,  145,  261,  792,  131,    5,    4,   72,   35,  148,    3,   15, 
         176,  485,  126,  142,    7,    9,   19,  977,   62,  142,   15,    1,  648,  237,    4,  369, 
          30,  134,    6,   15,    1,  644,  955,    0,    0,  925,  124,  171,    0,    0,  544,   28, 
         482,  482,  482,  131,  952,  380,  984,   76,   31,   72,   19,   68,  984,  316,  920,  936, 
         580,  593,    6,  845,  444,  738,  127,  577,   12,  652,   59,  644,  920,  936,  580,  389, 
           6,  648,   12,  971,  851,  577,   12,  772,  644,   12,   31,    8,  899,    4,  920,  936, 
         777,  184,  867,   78,  230,  444,  174,  697,   12,    0,   74,   84,   92,  111,  470,  714, 
         118,  125,  333,  837,  828,  140,  146,  152,  158,  164,  170,  178,  187,  194,  200,  204, 
         570,  209,  224,  231,  237,  243,  249,  257,  265,  636,  270,  811,  276,  292,  301,  306, 
         309,  318,  327,  355,  340,  346,  363,  369,  380,  386,  392,  282,  401,  409,   50,   69, 
         403,  375,  414,  552,  420,  422,  544,  428,  441,   79,  816,  456,  675,  476,  487,   97, 
         492,  578,  521,  508,  608,  526,  448,  287,  558,  594,  599,  604,  434,  613,  617,  621, 
         625,  631,  648,  823,  658,  664,  670,  688,  697,  680,  705,  218,  533,  642,  720,  726, 
         782,  732,  744,  751,  794,  788,  738,  776,  758,  800,  588,  764,  808,  107,   42,    0, 
         200,  396,  292,  265,  231,  536,  658,  194,  670,  675,  487,  295,  845,  992,  840,  158, 
        1004,  952,  572,  856,    8,  920,  892,  936,  992,   78,  624, 1016,  992,  133,  181,  992, 
        1023,  672,  176,  702,    0,   29,   96,  112,  992,  762,   23,   78,  672,  860,  758,  928, 
         614,  566,  630,   27,  550,  992,  502,   27,   78,   43,   74,  618,   86,  980,  980,  992, 
          74,   84,   92,  111,  776,  800,  758,  621,  625,   50,   69,   79,   97,  492,  476,  448, 
         422,  107,  664,   42,  570,  327,  428,  714,  355,  648,  636,  642,  152,  125,  170,  811, 
         470,  118,  340,  732,  794,  544,  744,  782,  375,  380,  270,  526,  409,  403,  599,  816, 
         243,  764,  578,  249,  608,  594,  552,  257,  788,  738,  823,  751,  441,  434,  178,  224, 
         276,  287,  282,  318,  533,  604,  187,  209,  146,  508,  237,  837,  828,  456,  521,  333, 
         558,  218,  688,  697,  680,  705,  414,  301,  726,  631,  164,  140,  369,  613,  309,  720, 
         999,  509,  188,  750,  961,    2,  661,  190,  617,  204,  392,  363,  386,  346,  803, 1008, 
         413,   88,  348,   14,  174,  752,  174,  622,  624,  980,  916,  971,  992,  933,   80,  323, 
         306, 1004,   78,  624,  888,   60,  262,    2,  992,  796,  746,  864,  572, 1003,  588,  420, 
         401, 1006,  110,  408,  174,  865,   80,  174,  672,  766,  928,  574,   51,  638,  992,    0, 
         808,    0,  981,  136,   24,  949,   80,  953,    2,  949,   80,  949,   80,   78,  624,   56, 
         174,  120,   40,  184,  104,  248,  168,  174,  232,  992,  672,   78,  622,  608,  494,  992, 
         327,  369,  270,  387,  321,  320,  322,  323,  328,  368,  270,  256,  376,  326,  325,  359, 
         352,  373,  480,    0,   23,   20,   17,   16,  339,  332,  271,    0,  424,  390,  412,  370, 
         338,  345,  401,   28,   24,   21,   18,   26,  337,  348,  463,  406,  425,  334,  413,  374, 
         342,  346,  400,   27,   25,   22,   19,  261,  343,  349,  464,  389,  428,  335,  414,  408, 
         336,  347,  264,    0,  268,  268,  268,    0,  341,  350,  263,  375,  268,  268,  268,    0, 
          65,   70,  270,   78,   81,   85,   89,   58,   97,  126,  270,   94,   45,   43,   42,   47, 
          66,   71,   75,    0,   82,   86,   90,   32,   98,   37,  127,    0,   55,   52,   49,   48, 
          67,   72,   76,   79,   83,   87,   61,   44,   99,   29,  410,   13,   56,   53,   50,   46, 
          68,   73,   77,   80,   84,   88,   63,  261,  100,   60,  411,   36,   57,   54,   51,  382, 
          69,   74,  264,    0,  268,  268,  268,    0,  101,   62,  519,  391,  268,  268,  268,  904, 
         238,  865,   80,   27,  986,  550,  758, 1007,  285,  100,  408,  916,   23,  980,   74,  250, 
         238,  344,  174,  270,  752,  668,   74,  604,  746,   39,  284,   80,  604,   14,  266,   74, 
        1006, 1006, 1006,  860,  550,  550,  358,  834,   31, 1018,    6,  738,   71,  764,   70,  550, 
         738,   31,  764,   70,  908,   19,  446,  112,  408,   29,   96,  344,  270,   56,  166,  262, 
         986,  614,   31,  762,  999,   70,  538,  433,   96,  752,  648,  408,  174,  908,   83,  133, 
          80,  672,  176,  750,  467,  574,  283,  443,  133,   80,  652,  151,  672,  176,  574,  379, 
         203,  133,   80,  750,  171,  867,   14,  176,  123,  248,  865,   80,  112,  176,  750,   83, 
         867,   14,  176,  203,  184,  174,  248,  878,  183,  716,  111,   78,  624,  952,  984,   76, 
          63,  984,  652,   39,  429,  112,   98,  961,    2,  184,  174,  248,  878,  871,  608,  716, 
          67,  321,  164,  997,  168,  189,  140,  899,   78,  624,  952,  984,   76,  935,  984,  652, 
         831,  429,  112,  100,  795,  206,  944,  750,  655,  811,  238,  880,   43,  206,  686,    0, 
         944,  936,  174,  344,  369,   28,  408,  174,  992,  176,  421,   88,  176,  174,   78,  624, 
         888,  444,   70,  518,   60,  872,  992,  888,  444,  174,  304,    5,  608,  518,   25,  114, 
         238,   56,  672,  558,  622,  766,   67,  574,   47,   56,   94,  574,   83,  638,  758,   27, 
          86,  630,  860,  738,   23,   78,  608,  238,  270,  752,   56,  878,   51,  588,  897,   11, 
         201,   10,  206,  752,  174,  992,  206,  638,  766,  187,  161,   24,  716,  864,  952,  856, 
          76,  864,  652,  928,  264,   65,  176,  952,  828,  856,  776,  328,  920,  764,  936,  992, 
          70,  624,  860,  160,  980,  980,  852,  815,  206,   88,  224,  412,  722,   81,  181,  931, 
         920,  572,  920,  764,  856,  952,   60,  984,  908,   19,  558,  780,   27,  558,  558,  444, 
         755,  885,   88,  304,    5,  885,   88,  304,    8,  885,   88,  304,    7,  856,  952,  700, 
         984,  780,  928,  964,  728,  856,   78,  304,  255,  984,  444,  270,  124,  672,  702,  608, 
        1009,   88,   91,  101,  115,  135,  161,  201,  267,  319,  399,  533,  432,  538,  816,  166, 
         638,  103,  638,  119,  638,  143,  286,  728,  446, 1019,  422,  987,  992,  728,  422, 1011, 
         992,  728,    0,  422, 1003,  992,  728,    0,    0,  422,  995,  992,  169,   92,  920,  444, 
         365,   30,  169,   92,  904,  971,  169,   92,  776,  939,  952,   60,  856,  900,  772,  992, 
         260,   78,  624,  888,   60,   90,  624,  174,   56,  238,  174,  270,  752,   56,  878,  864, 
         238,  268,   19,   78,  752,  366,  174,  891,  469,   92,  852,   43,  540,   82,  752,  992, 
          78,  752,  212,  864,  174,  624,   56,  988,  988,  988,  988,  915,  469,   92,  852,   75, 
         572,  732,   80,   16,  240,  624,  240,  827,  212,  967,  174,  624,   56,  988,  170,  988, 
         988,  892,  404,  995,  875,  304,    8,  624,  174,  224,  732,  160,  348,   56,   82,   28, 
         430,  750,  111,  174,  270,  624,   56,  980,  916,  955,  860,  754,  864,  220,  992,  924, 
         980,  980,  754, 1003,  992,  584,  166,  112,  645,   20,  344,  193,   92,   78,  624,  142, 
         888,   60,  454,  176,  454,  127,  264,  206,  174,  344,  590,   60,  230,  444,  238,  888, 
          90,  634,  174,  195,  408,  518,   55,  588,    9,  131,  584,  992,  888,  518,  444,  238, 
          90,  570,  174,  344,  888,  230,   43,  444,  538,  238,  752,  238,  174,  268,   51,  774, 
          51,  174,   46,   99,  870,  995,  174,  624,  250,  444,  538,   60,  230,   56,  238,   60, 
         624,  870,  815,  238,  752,  408,  238,  321,  164,  204,   23,  294,  110,  888,  518,   60, 
         518,  316,  518,   60,  872,  110,  580,   53,  190,  952,  856,   72,  920,  936,  992,    0, 
          78,   27,   78,  702,  860,   80,   27,   46,  122,  472,  408,   70,   62,   94,  472,  796, 
         980,  374,  566,  852,  995,  238,  750,  363,  472,  110,  750,  331,  806,  135,  472,  110, 
         806,  991,  174,  472,  782,   35,  472,  174,   43,  472,  174,  472,  110,  414,  862,   91, 
         654,  286,  806,   59,  472,  764,  472,  110,  422,  110,  806,   75,  358,  974,  190,  286, 
         980,  724,  963,   78,  174,  408,  238,  302,  630,  630,  630,    0,  203,   46,  122,  472, 
         408,   70,   62,   94,  472,  518,  606,   19,  670,   14,  472,  732,  988,  910,   19,  302, 
         610, 1011,  852,  971,  408,  174,  472,  408,  766,   27,  358,  974,  174,  860,  842,  191, 
         238,  174,  860,  270,  486,  107,  570,   91,  198,  550,  546,  222,  110,  762,  864,   78, 
          30,  992,  198,  963,  110,  867,  834,  847,  614, 1002,  995,   46,  250,  174,   78,  472, 
          78,  860,   80,  238,  174,  472,  174,   51,   46,  122,  472,  408,   70,   62,  762,  291, 
         472,  582,  606,   19,  670,  472,   94,  174,  110,  814,   43,  472, 1006,  614,  472,  860, 
          78,   19,  546,  398, 1011,  302, 1006,  980,  724,  979,  174,  408,  449,   98,   46,  250, 
         174,  862,   27,  181,  162,   62,  206,  110,  494,  494,  526,  238,   90,  270,  494,  486, 
          19,  698,  334,  924,  834,   23,  942,  910,   78,  110,  732,  336,  974,   83,  546,  462, 
        1011,  334, 1006,  916,  457,   99,  980,  970,  955,  422,   59,  707,  766,  695,  758,  679, 
         270,  142,   28, 1006,  906,  860,  842,  919,  358,  774,   27,  566,  992,   78,  546,  974, 
         574,  238,  706,   27,  938,  550,   14,  450,   35, 1006,  302, 1019,  478,   51,  906,  366, 
         550,  302, 1019,  106,  610,  875,  638,  859, 1006,  134,   90,   94,  298,  334,  186,  992, 
          78,  624,  158,  206,  616,  696,  166,  262,  680,  992,  126,  632,  238,  616,  696,  166, 
         126,  955,   78,  624,  632,  254,  472,  696,  222,  472,  992,  285,  100,  140,  437,   98, 
         408,  916,   31,  980,   74,  457,   98,   46,  250,  174,  732,  206,  472,  110,  206,  758, 
         864,  550,  742,   59,  614, 1006,   30,  980,  846,  975,  614,  992,  374,  762,   59,  566, 
         894,   19,   72,  582,   35,  438,  174,  147,   46,  240,  190,  240,   30,    6,  250,  398, 
        1019,  302, 1006,  614,  987,  910,  176,  437,   96,   76,  928,  762,  928,  270,  248,   29, 
          98,   14,  617,  100,  238,  176,  317,   96,  597,  100,  617,   98,  270,  597,  100,  309, 
          96,  617,  100,  629,   98,   78,  860,  550,  592,  992,   78,  472,  645,  100,  494,  974, 
         992,  860,   78,  464,  528,  336,  208,  592,  528,   80,  400,  208,  208,  592,  464,  336, 
         860,  992,  762,  928,  270,  142,  550,  550,  262,  860,  326,   71,  980,  916,   27,  206, 
         992,  614,  979,   78,  218,  140,  147,  988,  724,   35,  925,  100,   43,  988,  925,  100, 
         980,  980,  925,  100,  270,  206,  405,   98,   14,  917,  100,  988,  724,   23,  988,  917, 
         100, 1006,  334,  238,  915,  970,  522,  266,  970,  490,  490,  586,  140,   51,   14,  262, 
         526,   70,  992,  330,  970,  746, 1007,  992,  702,  110,  142,  472,  408,  910,  846,   39, 
         408,  270,  992,  550,  971,  860,  354,  110,  677,   98,   46,  250,  174,    4,  862,   19, 
           8,   30,   26,  110,  206,  486,  115,  206,  862,  127,  732,  980,  148,  389,  107,  550, 
         987,  757,  104,  419,  697,  104,  348,   51,  110,  358,  942,  819,  570,  398, 1011,  302, 
        1006,  614,   83,  156,  738,   43,  610,  738,   79,  546,  860,  291,  174, 1018,  174,  738, 
         875,   78,  860,  618,  270,  540,   80,   12,   19,  678,  110,  270,   76,   27,    9,   96, 
         652,   27,  702,  286,  529,   98,  546,  398, 1011,  302,  340,   63, 1006,  614,  980,  238, 
         523,  238,   76,   43,  553,  104,  174,  110,  732,  400,  156,  762,  411,  988,  738,   51, 
         610,  142,  472,  408,  131,  550,  910,  638,  923,  974,  974,  974,  354,  110,  270,   12, 
         569,   97,  595,  942,  638, 1011,  302,  382,  408,  811,  472,  408,  142,  238,  494,  494, 
         526,  110,  974,  750,   39,  408,  174,  992,  358,  971,  654,  472,  550,  661,   98,  110, 
          90,   94,  270,   12,   27,  993,  100,   76,   31,    1,   96,  321,  106,  238,  860,  144, 
         208,   16,  144,  336,  528,  336,   16,  592,  144,  592,  592,  272,  267,   78,  852,  151, 
         634,  272,  570,  212,  231,  596,  319,  276,  399,  660,  463,  340,  511,  924,  208,  348, 
         107,  400,  592,  208,   80,  272,  464,   80,  528,   16,  336,  400,  860,  238,  992,    0, 
         208,   80,   16,   80,  464,  592,  528,   16,  272,  208,  208,  412,  907,  284,  208,  208, 
          16,  528,  336,  208,   80,  400,  528,  220,  811,  348,  208,  208,  208,   16,  528,  208, 
         336,  604,  731,   92,  208,  208,  208,  208,   80,  284,  667,  540,  208,  208,  208,  668, 
         619,   46,  250,  174,  137,  100,  184,  865,   80,  270,  248,  862,  187,    6,  186,  758, 
          51,  781,   98,  742, 1003,  614, 1006,  858,  991,  742,   79,  190,  286,  510,  510,  542, 
         766,   19,  648,  184,   94,   46,  250,  174,  776,  730,  119,  209,  100,  762,  795,  408, 
         766,  775,   46,  529,   98,   46,  250,  174,   62,  862,  703,  730,  683,  166,  262,  742, 
         131,  326,   27,  678,    8,   14,   94,   90,  860,  394,  610,  546,  142,  472,  408,  395, 
         860,  206,  610,  174,  846,  845,  110,  834,   39,  614, 1006,  995,  472,  677,   96,  139, 
           1,   96,  691,   46,  250,  270,  174,  270,  550,  486,  947,  862,   87,  174,  997,  100, 
         860,   78,  166,  270,  110,   59,    8,  971,  340,  503,  980,  574,  550,  987,  627,  910, 
         638, 1011,  408,  302,  446,  563,  574,  110, 1006,  980,  148,  523,  174,  142, 1002, 1002, 
        1002,  174,  924,  464,  646,  710,  483,  348,  910,  238,  757,  104,  933,  108,  762,  227, 
         724,  955,   46,  924,  130,  302,  910,  693,  104,   12,   55,  110,  398,  110,  302,  110, 
          28,  933,  108,  762,   59,  910,  987,  238,  219,  910,   35,  862, 1007,  614,   94,   12, 
          27,  702,    0,  437,   96,  780,  203,  209,  100,  329,   96,  408,  766,   53,  106,  422, 
         238,  987,  910,  553,  104,  110,  348,  539,  302,  610, 1011,   66,  550,  988,  992,  140, 
         928,   78,  472,  697,  104,  238,  629,   98,   14,  697,  104,  176,  317,   96,  747,    0, 
           0,    0,    0,  176,    9,   70,  584,   22,  374,  790,  897,   11,  624,  449,   90,  257, 
          12,   16,    8,    1,   32,    4,    1,   20,    1,  260,    1,   20,    1,   32,    5,   18, 
          18,   15,   18,  269,    5,   13,   15,   18,   25,   32,   12,   15,   19,   20,  270,   15, 
          14,    5,   24,    9,   19,   20,    5,   14,   20,  270,   21,   12,   12,  272,   18,    9, 
          22,    1,   20,    5,  271,   21,   20,   32,   15,    6,   32,   18,    1,   14,    7,    5, 
         272,    1,    3,   11,    9,   14,    7,  276,   18,   25,   32,    1,    7,    1,    9,   14, 
         281,    5,   19,  270,   15,  274,    1,   13,  274,   15,   13,  264,  432,  608,  816,  570, 
         368,  444,  348,   80,  784,  270,  961,  176,  174,  816,  634,  262,   86,  936,  854,  979, 
         329,   36,  268,  928,  909,  444,  497,   14,  801,  112,  184,  240,  176,  270,   76,   35, 
         957,  112,   27,  949,  112,  873,  112,  909,  112,  176,  270,  309,   96,  873,  112,   76, 
          35,  953,  112,   27,  945,  112,  897,  112,   70,  624,  248,   76,   31,   72,  747,  270, 
         184,  309,   96,  873,  112,  941,  112,  897,  112,   14,  354,  873,  112,  937,  112,  909, 
         112,  240,   78,  624,  248,  296,   13,  114,  413,   88,  348,  238,  865,   80,  608,  238, 
         614,  624,  238,   56,  980,  916,  947,   78,  624,  275,  140,  928,  190,  702,  190,  992, 
          37,   96,   27,   29,   96,  165,   80,  752,  860,  992,  980,  980,  980,  980,  980,  608, 
          78,  624,  888,  444,  550,  988,  724, 1003,  614,  624,   56,  672,  860,  992,  801,  112, 
         949,  112,   29,  116,  240,  957,  112,  270,  937,  112,  238,   78,  624,  238,  609,   98, 
         132,  801,  112,  945,  112,  270,  937,  112,  309,   96,  129,  100,  140,   39,  949,  112, 
          27,  957,  112,  270,  309,   96,  702,  190,  201,  100,   49,   96,  937,  112,  617,   96, 
         129,  100,  937,  112,   46,  250,  270,    9,   96,  201,  100,  589,   96,  766,  649,    3, 
         773,   96,  140,  864,  240,  136,  953,  112,  619,  176,  762,  307,  766,   35,  648,  904, 
          94,  240,  270,  309,   96,  137,  100,  184,  270,  309,   96,  209,  100,   49,   96,  773, 
          96,  240,  270,  184,  174,  609,   96,  762,  223,   14,  203,  908,   31,  904,  992,  900, 
         992,  174,  648,  766,   19,  328,   94,  240,  176,  762,  928,   14,  491,  429,  116,  995, 
          46,  270,  122,  766,   75,  328,  524,   51,  908,   35,  900,  648,  324,  860,  166,  262, 
         486,  945,  119,  838,  143,  206,  718,  803,  860,  610,  750,   87,  780,  775,  645,  100, 
          14,  422,  174,   61,  122,  780,  781,   99,  569,   96,  429,  116,  110,  206,  860,   90, 
          94,  550,  742,   67,  574,  980,  340,  979,  238,   61,  122,  472,   78,  574,  974,  107, 
         174,  472,  546,  286,  472,  942,  942,  446, 1003,   30,  302,  174,  142,  462,  915,  472, 
         574,  472,  110, 1006,  980,  340,  947,  238,  701,   96,  110,  472,   70,  668,  238,  225, 
         120,  238,   19,  302,  610, 1011,  910,   66,  762,  283,  988,  923,  780,  227,  137,  100, 
           1,   96,  169,  100,    9,   96,  209,  100,  329,   96,   30,  773,   96,  176,   94,  472, 
         408,   70,  589,   96,  166,  262,  486,  673,  118,  689,  118,  988,  614,  852, 1003,   94, 
         437,   96,  908,   59,  702,  190,  617,  100,   49,   96,  652,   43,  617,  100,   49,   96, 
          76,  135,  617,  100,  358,  358,    0,  629,   96,  140,   63,   78,  860,  614,  592,  317, 
          96,  332,   19,  702,  524,  864,  240,  992,   78,  622,   94,  852,  111,  404,  239,  212, 
         295,  596,  335,  276,  359,  924,  464,  668,  992,  220,  400,  400,  528,  400,  336,  144, 
         272,  592,   80,   80,  400,  860,  992,  400,  916, 1011,  867,  284,  349,  120,  924,  336, 
          92,  528,  412,  992,  348,  349,  120,  924,  592,  220,  992,   92,  349,  120,  604,  992, 
         540,  349,  120,  284,  992,  520,  776,  174,   14,   46,  186,  766,   67,  648,  780,   27, 
         908,   19,  328,   94,  238,   76,  837,  123,  140,   43,  174,  270,  974,  462,   78,  860, 
         272,  336,  238,  614,  758,   47,  614,   27,  550,  910,  238,  472,  408,  494,  494,  494, 
         974,  238,  758,  159,  398, 1019,  302, 1006,  614,  987,   78,  238,  408,  494,   76,   27, 
         910,  974,  238,  398,   91,  302,  238,  408,  238,   76,  267,  742,  247, 1006,  235,  908, 
          71,  904,  332,   31,  328,  883,  324,  867,  900,  780,  963,  652,   27,  644,  811,  648, 
         795,  645,  100,  579,  110,  398,    0,  429,  116,   59,  550,  758,   39,  398,  947,  302, 
         614,    0,  437,   96,   76,   95,  408,  494,  614,    0,  617,   96,  617,  100,  329,   96, 
         472,  174,  270,  550,   59,  110, 1006,   59,  980,  340,  439,  550,  995,  110,   78,  238, 
         225,  120,  238,   19,  574,  398, 1011,  302,  980,  974, 1006,  340,  923,  472,  910,  910, 
          78,  860,   80,  472,  924,  400,  400,   91,  906,  906,  446, 1003,   30,  472,  174,  590, 
         302,  472,  142,  286,  610,  939,  174, 1018,  174,  762,  267,  638,  614,   30,  910,  923, 
         408,  524,  335,  908,  315,  569,   96,  291,  176,  472,  408,   70,  589,   96,  240,  209, 
         100,  329,   96,  908,   19,  240,  652,   19,  702,  240,  267,   94,  472,  174,  408,  430, 
         524,   31,  908,   31,  646,  110,  730,  195,  472,  677,   96,  780,  123,  137,  100,  209, 
         100,  329,   96,    1,   96,  773,   96,  524,  647,  569,   96,  332,  928,  702,  992,   78, 
         860,  618,   86,  270,  142,  780,  928,  803,    0,  237,  100,  762,  781,   99,  176,   76, 
         415,  270,   30,   78,  860,  614,  208,   29,   96,   78,   80,   16,  464,  208,  464,  272, 
          80,  528,  144,  272,  924,  592,  617,   96,  758,  781,   98,  224,  284,  160,  924,  110, 
          19,  910,  550, 1011,   78,  174,  494,  494,  494, 1006,  764,  160,  162,  224,  974,  980, 
         852,  939,  275,  924,   66,  742,  781,   99,  176,  546,   31,  986, 1003,  174,  418,   78, 
          46,  860,  528,  860,  238,  802,   39,  781,   98,  558,  418, 1011,  422,   55,  494,  494, 
         494, 1018,  923,  174,  176,   74,  796,   80,  144,  437,   98,  176,  262,   78,  304,  341, 
         892,  518,  892,  816,  992,  329,   36,  952,  572,  984,  908,   31,  904,   19,  900,  984, 
         892,  936,  992,  304,   45,  924,   88,  160,   81,  182,  408,  988,  208,  971,    6,  192, 
        
         580,   19,  584,  429,  112,   86,  569,   12,   81,  132,   78,  344,   68,  648,  929,  128, 
         917,  188,  752,  179,  213,  136,  138,  574,   35,  742,  983,  171,  170,  266,  112,  845, 
         164,  638,  892,  897,  188,  141,  140,  176,  170,  313,  136,  883,  777,   80,   78,   91, 
         268,  991,  408,  746,   45,  190,  266,  252,  845,  164,  857,  164,  170,  266,  344,  809, 
         164,  138,  321,  164,  204,   87,  408,  774,   71,  870,   47,  770,   39,  866,   19,   10, 
         174,  252,  202,  112,  260,  176,  266,  138,  176,  202,  112,  741,  164,  892,  738,   31, 
         758,  947,  610,  191,  610,  171,  502,   43,  502,   27,  758,  127,  268,   91,  408,  266, 
          70,  141,  140,  857,  164,  408,  170,  344,  264,   19,  260,  176,  266,  124,  774,  271, 
         870,   47,  770,  239,  866,  219, 1013,  168,  176,  170,  112,  741,  164,  234,  408,  624, 
         796,  161,  140,  408,  610,   35,  610,  610,  622,  610,  344,  176,  874,  887,  341,  130, 
          70,  252,  112,  138,  408,  266,  809,  164,  189,  140,  106,  731,   32,  176,  624,   56, 
         924,   88,  408,  624,  270,   56,  142,  910,  796,  438,   63,  438,  988,  988,  987,  258, 
         123,   74,  752,   28,  106,  272,   28,  770,  955,  166,  614,  624,  266,   78,  752,  408, 
         124,  170,  617,  140,  624,   56,  924,  152,  752,   70,  624,  888,  166,  872,   46,  870, 
         781,  186,  614,  624,  238,  752,  238,  963,   70,  624,  888,   28,  272,  624,   28,  266, 
          56,  992,  313,  136,  574,   55,  510,  510,  510,  689,  131,  408,  266,  124,  170,  617, 
         140,  252,  845,  164,  170,  344,  176,  266,  845,  164,  170,  266,  112,  741,  164,  892, 
         546,  477,  175,  992,  888,  230,   78,  304,  192,  344,  112,  131,  624,   56,  574,  147, 
         796,  746,   39,  380,  746,   35,  369,  132,   27,  341,  132,  198,  262,  176,  870,  879, 
         992,  638,  750,  928,  254,  220,   88,  176,  152,  112,  796,  176,  252,  618,  879,  124, 
         112,  341,  132,  734,  377,  133,  939,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
           0,    0,    0,    0,    0,  176,  624,  558,  112,   56,   14,   59,  341,  132,  408,  624, 
         558,  344,  174,  752,  992,  632,  344,  750,  139,  789,  152,  750,  897,   10,  588, 1007, 
         524,   39,  981,  136,  103,   28,  433,   24,   43,  204,  963,  425,   24,  174,  444,  816, 
         630,  630,  630,   39,  981,  136,   67,  634,  250,  645,   20,  262,  218,  282,  816,  774, 
           9,  131,  614,  230,   70,  624,  888,  624,  614,  444,  250,   56,  984,  132,  984,  752, 
         186,  570,  816,  796,  610,  258,  892,  162,  572,   14,  570,  816,  266,  638,   39, 1006, 
        1006,  971,  238,   60,  624,  614,  238,  174,  752,  238,  444,  614,   63,  238,  174,  732, 
         400,  796,  827,   60,  550,  262,   70,  624,  888,  166,  872,   28,    2,  196,  189,  140, 
         777,  184,  797,    2,  952,   70,  572,  856,  324,  644,  176,  992,  354,  857,  166,  366, 
         992,  196,   97,  164,  202,  984,  324,  984,  133,  164,  316,  266,  493,   26,  204,  928, 
         981,  136,  106,  614,  928,  140,  743,   70,  992,    0,    0,    0,    0,    0,    0,    0, 
          56,  363,   56,  291,   56,  259,   56,  227,   56,  195,   56,  163,   56,  252,  992,    0, 
          56,  992,   56,  147,   56,  115,   56,   83,   56,   51,   56,  915,   56,  892,  992,  316, 
         992,  380,  992,  124,  992,  572,  992,  134,  234,  614,  624,   56,  202,  992,  134,  230, 
         614,  624,   56,  198,  843,   66,  490,  490,  490,  546,  482,  486,   31,  966,   27,  966, 
         566,  522,   27,  550,   27,  610,  610,  266,  624,  124,  304,  544,  252,  480,  170,  963, 
         380,  984,  780,  745,   47,  885,  136,  889,  160,  389,   20,   12,  461,    7,  793,    2, 
         380,  984,  780,  721,   47,  885,  136,  321,  164, 1016,   12,  131,  742,  989,  169,  101, 
          80,  332,   19,   70,  550,   19,  614, 1000,  221,  140,  763,  742,   31,  550, 1000,  357, 
          20,  588,  793,   56,  101,   80,  550, 1000,  997,   92,  117,    6,  632,  344,  750,  135, 
         204,  287,  321,  164,  161,  164,  901,  132,  973,  168,  136,   78,  614,  584,  267,  789, 
         152,   28,  750,   27,  524,  891,  897,   10,  174,  614,  399,  132,   12,  371,   27,  136, 
          78,  112,  844,  327,  204,  713,  143,  321,  164, 1016,  973,  132, 1000,  580,  176,  324, 
         112,   25,  140,  332,   39,  176,  614,  971,  149,  164,  124,  170,  252,   97,  164,  124, 
         266,  588,  681,  167,  101,   80,  742,   35,  408,  941,  160,  797,    2,  837,  444,  529, 
          12,  369,   28,  557,  168,  844,  943,  992,  569,   12,  264,  608,  700,  856,  524,  928, 
         516,  920,  700,  936,  827,  929,  136,  432,  816,  453,  112,  716,   31,   76,   27,  889, 
         160,  669,   12,  557,  168,  891,  170,  266,  344,   72,  648, 1013,  168,  408,  170,  344, 
          51,   78,  857,  164,  141,  140,  408,  874,  975,  992,  170,  138,  624,  266,  124,  304, 
         643,  252,  480,  174,  796,  138,  624,  270,  124,  304,  640,  947,  797,  164,   75,  716, 
          63,   78,  624, 1016,   70,  614, 1000,   70,  624,  824,  170,  266,  204,   87,  482,   19, 
         546,  482,   19,  546,  482,   19,  546,  808,  992,   76,  969,  130,  857,  164,  157,  164, 
         170,  266,  809,  164,  170,  344,  313,  136,  574,   95,  328,  140,   51,  638,  510,  510, 
         510,  227,  432,  992,  408,  238,  845,  164,  741,  164,  796,  618,   79,  262,  998,   78, 
         624,  517,  188,  661,  188,  206,  344,   28,  266,  857,  164,  313,  136,  252,  238,  408, 
         124,  285,  136,  238,  124,  238,  106,  838,   23,   70,  566,  566,  518,   39,  630,  630, 
          19,  550,  106,  105,  140,  408,  266,  644, 1013,  170,  344,  842,   23,   74,  586,   35, 
         614,  610,  610,  486,  486,  486,  486,   19,  546,  970,  784,   28,  266,  408,  109,  140, 
         408,  992,  953,  132,  844,  529,  135,  174,  321,  164,  580, 1016,  742,   51,  997,  168, 
         332,   55,  584,  101,   80,  550, 1000,  221,  142,  816,  986,  986,  986,  494,  494,  992, 
         432,   43,  432,  570,  368,  634,  805,  140,  243,  432,   43,  432,  570,  368,  634,  805, 
         140,  163,  432,   43,  432,  570,  368,  634,  805,  140,   83,  432,   43,  432,  570,  368, 
         634,  805,  140,  570,  570,  570,  892,  494,  494,  480,  432,  368,  572,   70,  892,  480, 
         102,  444,  796,  570,  816,  630,  758,  999,  738,   63,  746,  963,  614,  874,  943,  259, 
         546,  546,  546,  546,  891,  924,  546,  159,  546,  847,  570,  570,  816,  796,  546,  807, 
          78,  588,  127,  584,  142,  425,   24,  110,  444,  715,  570,  816,  870,  687,  634,  634, 
          60,   28,  992,  324,  580,  134,  321,  164,  204,  575,  198,  444,   88,  332,   27,  845, 
         164,  741,  164,  892,  642,  482,  991,  482,  311,  482,  943,  482,   35,  477,  172,  915, 
         758,  899,  900,  630,  572,  174,  444,  924,  152,  278,   28,  870,  103,   60,  270,  809, 
         164,  908,  809,  165,   78,  624,  170,  992,   60,  270,  699,  857,  164,  675,  738,  999, 
         566,  199,  566,  967,  313,  136,  574,  935,  588,   47,  493,   24,  584,  547,  332,   59, 
         321,  164,  845,  164,  221,  140,   78,  624,  992,  741,  164,  904,  587,  893,  156,  408, 
         716,  191,   76,  175,  588,  155,  203,  860,   66,  750,  299,  270,   78,  624,  796,  842, 
          51,  170,  892,  910,  910,  979,  572,  344,  616,  789,  152,  750,  155,  524,   31,  196, 
         147,  588,  123,  140,  423,  344,  696,  742,  387,  952,  856,  408,  444,  816,  742,  331, 
         480,  200,   28,  266,  797,  164,  163,  893,  156,  644,   17,    0,  638,  766,  587,  909, 
           8,  262,  304,  100,  774,  155,  909,  144,   28,  266,  696,  742,  435,  138,   99,  106, 
         902,  902,  422,  324,  209,  144,  750,  864,  897,   10,   70,  624,  716,   47,  952,  856, 
          76,  131,  696,  266,  824,  170,  252,  270,  760,  252,  170,  744,  174,    9,   48,  171, 
         234,    1,   48,  777,   30,  772,  716,  127,   76,  111,  262,  408,  588,  909,  144,  780, 
         903,  266,  189,  140,  961,    2,  204,  307,  266,    2,  824,  444,  570,  816,  166,  182, 
         570,  816,  764,  486,   71,  824,  170,  458,  780,  843,  138,  571,  824,  330,  979,  776, 
         238,  321,  164,  829,  164,  829,  164,  170,  266,  853,  156,  238,  595,  268,   59,  234, 
         329,  164,  741,  164,  214,  742,  307,   66,  490,  490,  490,  546,  482,  486,  151,  966, 
         234,  941,   60,  472,  106,  652,  131,  326,  322,   83,  358,  408,  856,   70,  624,  587, 
         966,  566,  883,  418,  418,  947,  170,  610,  610,  781,  164,  899,  264,  941,   60,  644, 
         984,  262,  328,  913,  144,  266,  472,  870,   39,  770,   51,   27,  774,   27,  260,  170, 
         582,  578,   35,  614,  610,  610,  486,  486,  486,  486,   19,  546,  970,  230,  321,  164, 
         749,  164,  892,  198,  572,  250,  254,  141,  140,  857,  164,  206,  892,  141,  140,  741, 
         164,  984,  644,  268,   19,  648,  984,  141,  140,  408,  266,  373,  150,  537,    8,  854, 
         928,  138,   22,  204,  195,  838,  139,    2,  166,  856,  652,   59,  644,  920,  262,  824, 
         330,   75,  262,  824,  170,  458,   35,  893,  144,  266,   73,  150,  838,  187, 1002, 1002, 
         902,  902,  824,  482,  170,  482,   39,  781,  164,  907,  326,  546,  546,  322,   27,  358, 
         851,  418,  418,  827,  260,  893,  144,  344,  321,  164,  112,  408,  870,   39,  770,   51, 
          27,  774,   27,  264,  170,  781,  164,  854,  151,  998,  854,  127,  998,  906,  176,  170, 
         268,   19,  546,  490,  490,  490,  486,  572,  141,  140,  408,  805,  150,  540,  400,   60, 
         286,  408,  238,  106,  545,  176,    0,  796,  758,   27,  272,  796,  238,  234,  572,  746, 
          35,  446,   47,  891,  572,  746, 1011,  344,  132,  348,   78,  624,  336,  250,  218,  924, 
         816,   88,  570,  816,  742,   87,  348,  218,  546,  931,   80,  208,  976,  976,  136,  796, 
         570,  816,  140,  407,  230,  570,  816,  710,   31,  742,  867,  230,  270,  188,  322,  636, 
         166,  892,  202,  112,  444,  166,  502,  502,  502,  419,  570,  570,  270,  816,  828,  286, 
         632,  174,  638,  570,  570,  816,  874,  103,  638,  910,  910,  766,   47,  842,   47,  580, 
         483,  842,  919,  188,  611,   28,  262,  838,   31,   78,  992,  304,  991,  774,   71,  454, 
          60,    2,  522,  444,  261,  154,  166,  764,  970,  546,  796,  112,  444,  270,  408,  174, 
         634,  816,  746,  131,  260,  984,  652,   27,  644,  264,  984,  874,   63,  910,  910,  268, 
          79,  842,  887,  124,  140,   23,  828,  257,  154,  842,  975,  584,  176,  668,   16,  140, 
         159,  270,  572,  634,  634,  506,  506,  506,  986,  506,  506,  156,  152,  506,  506,  668, 
         656,   28,  170,  520,  992,  888,   28,  272,   28,  266,  624,   56,  572,  742,   53,  154, 
         213,  136,  574,  979,  636,  610,   88,  138,  202,  252,  202,  270,  845,  164,  857,  164, 
         408,  238,  110,  110,   28,  741,  164,  110,  796,  874,   87,  910,  910,  152,  610,   88, 
         738,   75,  842,  903,   28,  206,  124,  266,  188,  675,  842,  975,   70,  624,  206,  124, 
         516,  580,  992,  580,   28,  716,   31,   76,  315,  760,  270,  824,  170,  124,  746,  235, 
         200,  738,   71,  196,  490,  490,  490,  486,  111,  966,  808,  174,   74,  124,  744, 1016, 
          70,  614, 1000,  137,   10,  966,  566,  923,   78,  624,  584,  723,  708,  588,  928, 1016, 
          70, 1000,  204,   87,  149,  164,  316,  266,  493,   24,  580,   53,  190,  425,   24,  987, 
         566,  175,  819,  344,  566,  199,  566,  153,    3,  716,   31,   76,  931,  329,  164,  829, 
         164,   29,  180,  572,  574,  875,  408,  270,   70,  624,   17,   12,   27,  537,    8,  140, 
         864,  985,   28,  952,  329,   38,  630,  963,   33,    6,  632,  344,  750,  817,  158,  696, 
         170,  680,  789,  152,  750,  929,  146,  616,  696,  262,  509,  188,  750,   59,  696,  270, 
         776,  513,  172,   27,  661,  188,  696,  262, 1006, 1006,  632,  124,  238,  524,  255,  632, 
         174,  572,  238,   28,  845,  164,  857,  164,  705,  164,  110,  796,  874,  928,  110,   28, 
         344,  238,  141,  140,  796,  408,  746,  928,  174,   70,  624,  645,   82,  513,  172,   12, 
         864,   78,  202,  252,  170,  572,  638,  238,  797,  160,  750,   63,  624,  110,  645,   80, 
           9,  130,  624,  344,   56,  238,  752,  408,  550,  774,  963,  992,  142,  645,   80,  110, 
         776,  513,  174,  321,  164,  204,   47,   70,  970,  326,    2,  696,  170,  680,  992,  652, 
         927,    6,   28,  963,  304,   11,  262,  516,  952,  920,  936,  166,  828,  432,  764,   28, 
         272,  646,  444,  348,  546,   27,  124,  480,  816,  742,  979,  480,    0,    0,    0,    0, 
          56,  291,   56,  243,   56,  195,   56,  147,   56,   99,   56,   51,   56,  892,  202,  572, 
         179,  252,  202,  124,  147,  316,  202,  380,  115,  380,  202,  316,   83,  124,  202,  252, 
          51,  572,  202,  892,   19,  202,  752,   28,  992,  572,  234,  892,  291,  981,  136,   34, 
          56,  259,   56,  915,   56,  867,   56,  819,   56,  771,   56,  723,   56,  675,  627,    0, 
          56,  347,   56,  819,   56,  283,   56,  235,   56,  187,   56,  139,   56,  892,  234,  572, 
         235,  892,  194,  214,  572,  752,  170,  266,  622,  624,  796,  795,  252,  234,  124,  115, 
         316,  234,  380,   83,  380,  234,  316,   51,  124,  234,  252,   19,  234,  714,   71,  752, 
         408,  574,  174,   70,  624,  992,  785,  160,  750,  467,  165,  164,   97,  164,  124,  285, 
         136,  742,   19,  558,  105,  140,  408,  266,  828,  796,   35,  630,  988,  988,  630,  995, 
          78,  624,  888,  622,  872,  558,  624,  230,   56,  230,  614,  624,  230,  752,  230,  550, 
         870,  935,  230,  174,  752,   78,  170,  174,   56,  174,  752,  408,  624,   56,   74,  752, 
         408,  937,  166,  408,  266,   67,  809,  164,   70,  133,  164,  638,  344,  766,  967,  588, 
          19,  712,    9,  130,   78,   28,  624,  888,  622,  624,  262,   56,  750,   47,  304,  192, 
         774,  928,   78,  992,  204,  135,  149,  164,  316,  266,  177,  140,  577,  170,  557,  168, 
         614,  927,  742,  907, 1000,  321,  164,  204,  303,  161,  164,  472,  842,   39,  777,   80, 
          27,  809,  164,  749,  164,  892,  964,   72,   59,  252,  202,  174,  472,   81,  172,  472, 
         138,  174,  774,  951,  870,   47,  770,  919,  874,  899,  316,  969,  170,  444,  264,  816, 
         634,  630, 1007,   60,  638,  581,  170,  931,  344,  316,  266,  845,  164,  749,  164,  924, 
         976,  141,  140,  408,  992,  321,  164,  170,  472,  929,  128,  572,   27,  213,  136,  472, 
         774,   63,  870,  864,  770,   31,  866,  864,  124,  138,  202,  252,  472,  574,  103,  472, 
         316,  202,  380,  472,  836,  638,  510,  510,   19,  840,  742,  791,   10,   78,  472,  992, 
          78,  624,  824,   28,  204,   23,  482,  266,  992,   28,  174,  742,  189,  158,   90,  550, 
         143,  550,   59,  304,   29,  892,  580,  465,    2,  614,  614,  252,  264,  589,  168,  965, 
           2,  888,  272,   28,  266,  112,  313,  136,  742,   39,  777,   80,   59,  213,  136,  574, 
         111,  845,  164,  741,  164,  892,  738,   31,  758,  979,  176,  874,  219,  785,  160,  750, 
           9,  130,  156,  784,   28,  304,  288,  752,  176,  624,  614,  266,   56,  984,  132,  520, 
         984,  752,   78,  624,  888,  614,  872,  196,  177,  140,    1,  128,  189,  156,  961,    2, 
         204,   83,  174,  270,  444,  816,  992,  845,  164,  857,  164,  170,  266,  624,  124,  304, 
         545,  252,  480,  454,  450,  928,  187,   28,  204,  183,  354,  354,  354,  881,  134,  204, 
         143,   28,   35,  418,   55,  418,  418,   47,  418,  992,  418,  418,  418,  418,  418,  430, 
         992,  366,  992,   70,  924,   88,  837,  164,  174,  344,  624,  124,  924,  152,  230,  796, 
         304,  644,  252,  480,  713,  140,  142,  206,  860,   88,   30,  921,  164,  670,  510,   91, 
         574,  574,  187,  501,  168,  913,  164,  461,  168,  131,  510,  405,  170,  766,  503,  860, 
         546,   75,  252,  550,  796,  738,  463,  141,  140,  395,  546,  423,  260,  546,   23,  264, 
         909,  164,  304,   15,  268,   35,  913,  164,   83,  501,  168,  550,  913,  164,  909,  164, 
         461,  168,  321,  164,  857,  164,  157,  164,  617,  140,  124,  617,  140,  268,   99,  252, 
          97,  164,  266,  845,  164,  221,  140, 1016,   70, 1000,  965,    2,  510,  766,   55,  206, 
         220,  917,  164,  955,  860,  610,   67,  412,  738,  951,  144,  252,   93,  170,  610,  899, 
         412,  738,  879,  208,  955,  909,  164,  510,  766,  819,  252,  550,  796,  738,  783,  720, 
         797,  164,  851,  632,  750,  928,  913,  164,  632,  974,  974,  616,  963,  304,  240,  174, 
         344,  632,   35,  358,  974,  974,  750,  999,  408,  174,  992, 1016,  550,   31,  614,  992, 
         260,   78,  622,  160,   92,  224,  112,  204,  423,  149,  164,  268,   19,  316,   82,  472, 
         842,   67,   27,  213,  136,  574,   51,  742,  991,  777,   80,   51,  857,  164,  741,  164, 
         892,  964,   72,  138,  472,  270,  176,  202,  112,  174,  472,   81,  172,  472,  562,  174, 
         882,   75,  774,  943,  870,   47,  770,  911,  866,  891,  174,  227,  425,   24,   78,  170, 
         344,  426,  268,  321,  164,  176,  170,  472,  270,  324,   43,  997,  168,  332,   63,  370, 
         408,  786,   27,  778,  959,  174,  112,  124,  262,  101,   80,  160,   28,  844,  864,  166, 
        1000,  176,  266,  221,  140, 1016,  992,  964,   27,  964,  136,  204,   39,  741,  164,  259, 
         170,  444,  570,  816,  758, 1003,  570,  816,  630, 1007,  634,  630,  481,   27,  328,  140, 
         425,   26,  634,  955,  418,   75,  170,  610,  610,  614,  624,  266,   56,  892,  418,  892, 
         642,  482,  251,  546,  546,  928,  502,   43,  502,   27,  758,  847,  234,  202,  397,  172, 
         642,  482,   83,  546,  546,   59,  502,  939,  502,  923,  758,  907,  809,  164,  572,  202, 
         992,  482,  235,  738,  255,  566,  239,  566,  223,  652,  293,  143,  397,  172,  397,  172, 
         546,  311,  328,   76,  864,  809,  164,  809,  164,  140,  791,  313,  136,  493,   26,  482, 
         139,  397,  172,  418,   83,  170,  784,   28,  614,  624,  266,   56,  252,  992,  418,  892, 
         992,  482,   47,  758,  864,   81,  174,  630,  864,  234,  397,  172,  234,  630,  987,  515, 
           4,  888,   28,  272,  344,   28,  252,  202,  238,  304,  191,  550,  174,  472,  870,  363, 
         472,  174,  624,  112,   56,  574,  323,  638,  286,  796,  874,   35,  380,  874,  231,  842, 
         127,   28,  906,  906,  166,  182,  572,  202,    8,  380,  894,   19,  380,  752,   59,  780, 
          35,   74,  572,  947,  572,  472,   70,  624,  472,  992,  176,  643,  472,   19,  174,  252, 
         238,  112,  124,   28,  266,  313,  136,  742,  203,  213,  136,  574,  987,  252,  170,  270, 
         344,  845,  164,  741,  164,  138,  796,  218,  124,  266,  252,  874,  183,  842,   87,   70, 
          28,  218,  624,  124,  270,  176,  238,  627,  780,   51,   70,  110,  141,  140,  571,  408, 
           8,  547,   28,  408,  266,  124,  651,  304,   32,  262,  796, 1016,  874, 1011,  952,  992, 
         127,   97,   98,   99,  100,  101,    0,   96,    6,    4,    5,    1,   12,   29,  126,   13, 
          78, 1008,   92,  400,  304,  140,  828,  270,  741,  164,  796,  746,   87,  304,    5,   28, 
          66,  874,  951,  961,  176,  107,  572,  961,  176,  736,  299,  110,  304,    5,   28,   66, 
         874,  159,  158,  304,   31,  268,   35, 1000,  446,   55,  550,  446,   31, 1000, 1003,  736, 
         800,  222,  365,  186,  862,   39,  268,  881,  176,  329,   36,   28,  741,  164,  572,  142, 
         985,   28,  892,   86,  373,  176,  683,  304,  128,  163,  304,  192,  139,  262,   22,  304, 
          58,  870,  939,  304,   44,  870,  931,  304,   46,  870,  247,  304,   64,  262,  952,  984, 
         332,   95,  652,   79,  984,  732,  784,  286,  222,  894,   51,   83,  984, 1000,  304,   32, 
         734,   35,  126,  446,  126,  880, 1000,  992,   22,  304,   32,  774,  151,  304,   96,  774, 
         115,  166,  984,  324,  984,  262,  432,  816,  368,  166,  838,  928,    6,  795,   78,  348, 
         144,  784,   28,  816,  870,   51,  546,  995,  304,   58,  859,   60,   86,  566,  827,   14, 
         321,  164,  705,  164,  796,   66,  618,  864,  252,   92,  258,   29,  180,  142,  924,   88, 
         262,   22,   70,  624,  304,  127,  870,  901,   29,  206,  270,   28,  124,  614,  221,  143, 
         252,  270,   29,  180,  142,  924,   88,   70,  624,   81,  180,  883,  736,  800,  268,  864, 
         588,   63,  968,  972,   55,  584,  621,    0,  972,  864,  304,  896,  486,  614, 1019,  992, 
         304,   16,  624,  304,  253, 1008,  412,   74,  220,  144,  668,  144,   92,  144,  796,  144, 
         296,  296,  296,  992,  329,   36,  110,   28,  204,  741,  166,  366,  713,  166,  568,  796, 
         572,  746,  877,   89,  796,  568,  892,  270,  504,  892,  266,  174,  552,  440,  892,  266, 
         174,  488,  376,  892,  266,  174,  424,  174,  924,  152,  360,  992,  230,  293,   28,  230, 
          86,  262,  924,   88,  952,  380,  984,  772,  984,  316,  936,  502,  502,  303,  838,  135, 
         140,  231,   12,   35,  304,   11,  992,  652,   39,  304,  119,  992,  304,  135,  992,  304, 
          28,  870,   39,  304,   84,  992,  669,   88,   12,  713,   34,  393,  186,  132,  952,  920, 
         936,  299,  136,  952,  920,  936,   12,  423,  652,  171,  304,  127,  262,  924,  152,  742, 
         909,   38,  870,  175,  613,   32,  131,  952,  316,  984,  776,  984,  380,  936,  217,   32, 
         377,   36,  957,   32,  293,   36,  797,    2,   57,  180,  632,  766,   55,  254,  985,   28, 
         952,   27,  265,  184,   70,  152,  373,  176,  305,  184,  867,  652,   65,  187,  321,  164, 
          25,  140,   78,  624,  217,   32,  321,  164,   30,  142,  741,  164,  796,  746,   43,  110, 
         909,  164,   30,   70,  624,  524,   27,   41,  184,  224,  860,  160,  632,  672,  766,  123, 
         670,  608,  254,  222,  638,   91,  908,   75,  254,  304,   26,   49,  184,  947,  638,  608, 
         254,  224,  724,  343,  632,  546,  175,  532,   87,  610,  988,   80,   88,  980,  160,  921, 
         164,  787,  780,  119,  908,  195,  638,  183,  638,  167,  195,  788,  183,  916,  167,  780, 
         147,  796,  160,  304,   27,   49,  184,  632,  758,  595,   41,  184,  571,  160,  909,  164, 
         260,   43,  160,  909,  164,  264,  397,   20,  797,    2,  304,   28,  924,   88,  921,  166, 
         304,  127,  870,  915,  632,  838,  151,  638,  766,   47,  577,   12,  701,  138,  174,  141, 
         140,  809,  164,   70,  624,  174,  616,   99,  574,   35,  613,   32,  739,  174,  921,  164, 
         446,    0,  907,  286,  321,  164,  857,  164,  190,  286,  764,  796,  976,  141,  140,  382, 
         519,  547,  632,  286,  158,  985,   28,  862,  928,  446,  952,  995,  304,   31, 1000,  304, 
          32,  222,  638,  111,  286,  574,  862,   35, 1000,  446,  995,   70, 1008,  624,  616,  992, 
          94,  979,  952,  856,   12,  311,  316,  984,  904,  984,  380,  936,   70,  924,  152,  262, 
         304,  127,  870,  127,  376,  796,  746,   63,  732,  784,  254,  985,   28,   27,  265,  184, 
         609,  182,  901,   28,  732,  784,  254,  961,  176,  593,  182,  713,  140,  924,  152,  112, 
         321,  164,   30,  304,  241,  924,   88,  921,  164,  176,  924,   88,  921,  164,  174,  638, 
         616,   21,  186,   78,  624,  348,  784,   92,  976,  784,  270,  952,  944,  572,  262,  506, 
         506,  124,  326,  568,  444,  166,  262,  856,   60,  552,  992,  742,  279,   78,  112,  777, 
          80,  307,  580,  929,  128,  170,  112,    4,  266,  845,  164,  749,  164,  984,  780,   39, 
         260,  984,   51,  264,  772,  984,  141,  140,  176,  270,  313,  136,  742,  771,  213,  136, 
         574,  727,  170,  266,  112,  845,  164,  268,  235,    8,  749,  164,  892,  418,   75,  170, 
         610,  610,  614,  624,  266,   56,  892,  418,  892,  642,  482,  919,  482,  239,  482,  375, 
         482,  867,  477,  172,  843,  176,  742,  527,  624,   12,   75,  321,  164,   78,  624,  744, 
         808,  221,  140,  952,  856,  588,  928,  981,  136,   95,  482,  127,  738,  279,  566,   95, 
         566,   79,  857,  164,  741,  164,  892,  546,  727,  739,  397,  172,  523,  749,  164,  892, 
          86,  572,  141,  140,  741,  164,  796,   74,  238,  206,  141,  140,  206,  892,  867,  741, 
         164,  796,   74,  238,  206,  141,  140,  206,  892,  795,  166,  764,   88,  110,   29,  180, 
         540,  152,    1,   32,  195,  174,  444,  985,   28,   12,  115,  570,  570,  816,  262,  422, 
          60,  558,  238,  953,  188,  260,  981,   18,  845,   20,  521,   18,  985,   28,  953,  188, 
         206,   60,  262,   30,  929,   20,  952,  796,  976, 1000,  102,   30,  929,   20,  867,  422, 
        1006,  540,  272,  900,  528,  796,  578,   31,  258,  904,  156,   27,  988,  988,  438, 1003, 
         998,  790,   31,  988,  470,   78,  916,  864,  546,   19,  482,  438, 1011,  270, 1016,  908, 
          23,  696,  344,  944,  992,  750,   39,  408,  514,   35,  408,  174,  590,  752,  992,  206, 
         112,  152,  920,    1,   32,  123,   12,   63,  952,  856,  176,  174,  444,  480,  110,  845, 
         156,  206,  773,  146,  897,   10,   68,  260,  772,  524,   71,  837,  164,  741,  164,  857, 
         164,   43,  366,   45,  180,  366,  614,  230,  110,  985,   28,   76,  985,  176,  985,   18, 
         268,   35,  238,  344,  238,  260,  984,  524,   35,  264,  516,  776,  984,  992,  957,   28, 
          24,   18,   15,   13,  544,  992,    0,    0,    0,    0,    0,    0,    0,    0,    6,  237
          ,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,
           0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0           

    );
    signal raddr : integer range 0 to 16383 := 0;
begin

    Q <= std_logic_vector(to_unsigned(rom(raddr), 10 ));
    process(OutClock)
    begin
        if rising_edge(OutClock) then
            raddr <= to_integer(unsigned(Address));
        end if;
    end process;
    
end logic;
